VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dff_ram
  CLASS BLOCK ;
  FOREIGN dff_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.000 BY 2000.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 419.020 402.320 420.620 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 572.620 402.320 574.220 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 726.220 402.320 727.820 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 879.820 402.320 881.420 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1033.420 402.320 1035.020 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1187.020 402.320 1188.620 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1340.620 402.320 1342.220 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1494.220 402.320 1495.820 1599.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 421.710 1600.120 423.310 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 574.890 1600.120 576.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 728.070 1600.120 729.670 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 881.250 1600.120 882.850 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1034.430 1600.120 1036.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1187.610 1600.120 1189.210 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1340.790 1600.120 1342.390 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1493.970 1600.120 1495.570 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 415.720 402.320 417.320 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 569.320 402.320 570.920 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 722.920 402.320 724.520 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 876.520 402.320 878.120 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1030.120 402.320 1031.720 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1183.720 402.320 1185.320 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1337.320 402.320 1338.920 1599.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1490.920 402.320 1492.520 1599.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 418.410 1600.120 420.010 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 571.590 1600.120 573.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 724.770 1600.120 726.370 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 877.950 1600.120 879.550 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1031.130 1600.120 1032.730 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1184.310 1600.120 1185.910 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1337.490 1600.120 1339.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 399.960 1490.670 1600.120 1492.270 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 1996.000 982.470 2000.000 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END addr[1]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END clk
  PIN data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 646.040 2000.000 646.640 ;
    END
  END data[0]
  PIN data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 758.240 2000.000 758.840 ;
    END
  END data[10]
  PIN data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END data[11]
  PIN data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 1996.000 142.050 2000.000 ;
    END
  END data[12]
  PIN data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 1996.000 666.910 2000.000 ;
    END
  END data[13]
  PIN data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END data[14]
  PIN data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1996.000 824.690 2000.000 ;
    END
  END data[15]
  PIN data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END data[16]
  PIN data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 1996.000 1033.990 2000.000 ;
    END
  END data[17]
  PIN data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1989.040 4.000 1989.640 ;
    END
  END data[18]
  PIN data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END data[19]
  PIN data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1996.000 876.210 2000.000 ;
    END
  END data[1]
  PIN data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 1996.000 248.310 2000.000 ;
    END
  END data[20]
  PIN data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1421.240 2000.000 1421.840 ;
    END
  END data[21]
  PIN data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END data[22]
  PIN data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1876.840 4.000 1877.440 ;
    END
  END data[23]
  PIN data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1996.000 560.650 2000.000 ;
    END
  END data[24]
  PIN data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END data[25]
  PIN data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.240 4.000 1710.840 ;
    END
  END data[26]
  PIN data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1642.240 2000.000 1642.840 ;
    END
  END data[27]
  PIN data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1088.040 2000.000 1088.640 ;
    END
  END data[28]
  PIN data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END data[29]
  PIN data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 1996.000 1401.070 2000.000 ;
    END
  END data[2]
  PIN data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1972.040 2000.000 1972.640 ;
    END
  END data[30]
  PIN data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1587.840 2000.000 1588.440 ;
    END
  END data[31]
  PIN data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 812.640 2000.000 813.240 ;
    END
  END data[32]
  PIN data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END data[33]
  PIN data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.050 1996.000 1346.330 2000.000 ;
    END
  END data[34]
  PIN data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 1996.000 1661.890 2000.000 ;
    END
  END data[35]
  PIN data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data[36]
  PIN data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END data[37]
  PIN data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END data[38]
  PIN data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END data[39]
  PIN data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END data[3]
  PIN data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END data[40]
  PIN data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.240 4.000 1268.840 ;
    END
  END data[41]
  PIN data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 703.840 2000.000 704.440 ;
    END
  END data[42]
  PIN data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1254.640 2000.000 1255.240 ;
    END
  END data[43]
  PIN data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END data[44]
  PIN data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END data[45]
  PIN data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 979.240 2000.000 979.840 ;
    END
  END data[46]
  PIN data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 1996.000 1137.030 2000.000 ;
    END
  END data[47]
  PIN data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END data[48]
  PIN data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1996.000 927.730 2000.000 ;
    END
  END data[49]
  PIN data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 95.240 2000.000 95.840 ;
    END
  END data[4]
  PIN data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1696.640 2000.000 1697.240 ;
    END
  END data[50]
  PIN data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.950 1996.000 1974.230 2000.000 ;
    END
  END data[51]
  PIN data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 1996.000 718.430 2000.000 ;
    END
  END data[52]
  PIN data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 0.000 1516.990 4.000 ;
    END
  END data[53]
  PIN data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1475.640 2000.000 1476.240 ;
    END
  END data[54]
  PIN data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.130 1996.000 1713.410 2000.000 ;
    END
  END data[55]
  PIN data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 0.000 1465.470 4.000 ;
    END
  END data[56]
  PIN data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 1996.000 1922.710 2000.000 ;
    END
  END data[57]
  PIN data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1808.840 2000.000 1809.440 ;
    END
  END data[58]
  PIN data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1996.000 299.830 2000.000 ;
    END
  END data[59]
  PIN data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 37.440 2000.000 38.040 ;
    END
  END data[5]
  PIN data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END data[60]
  PIN data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END data[61]
  PIN data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END data[62]
  PIN data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 1996.000 196.790 2000.000 ;
    END
  END data[63]
  PIN data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END data[64]
  PIN data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1996.000 90.530 2000.000 ;
    END
  END data[65]
  PIN data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 1996.000 1294.810 2000.000 ;
    END
  END data[66]
  PIN data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END data[67]
  PIN data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 149.640 2000.000 150.240 ;
    END
  END data[68]
  PIN data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END data[69]
  PIN data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 479.440 2000.000 480.040 ;
    END
  END data[6]
  PIN data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.750 0.000 1620.030 4.000 ;
    END
  END data[70]
  PIN data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1917.640 2000.000 1918.240 ;
    END
  END data[71]
  PIN data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 591.640 2000.000 592.240 ;
    END
  END data[7]
  PIN data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END data[8]
  PIN data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END data[9]
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 1996.000 1555.630 2000.000 ;
    END
  END enb
  PIN r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 1996.000 509.130 2000.000 ;
    END
  END r_data[0]
  PIN r_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END r_data[10]
  PIN r_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1366.840 2000.000 1367.440 ;
    END
  END r_data[11]
  PIN r_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 370.640 2000.000 371.240 ;
    END
  END r_data[12]
  PIN r_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.090 1996.000 1610.370 2000.000 ;
    END
  END r_data[13]
  PIN r_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.010 1996.000 1243.290 2000.000 ;
    END
  END r_data[14]
  PIN r_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 1996.000 1819.670 2000.000 ;
    END
  END r_data[15]
  PIN r_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END r_data[16]
  PIN r_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END r_data[17]
  PIN r_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END r_data[18]
  PIN r_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END r_data[19]
  PIN r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1145.840 2000.000 1146.440 ;
    END
  END r_data[1]
  PIN r_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 867.040 2000.000 867.640 ;
    END
  END r_data[20]
  PIN r_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1996.000 773.170 2000.000 ;
    END
  END r_data[21]
  PIN r_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 1996.000 406.090 2000.000 ;
    END
  END r_data[22]
  PIN r_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 204.040 2000.000 204.640 ;
    END
  END r_data[23]
  PIN r_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END r_data[24]
  PIN r_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END r_data[25]
  PIN r_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END r_data[26]
  PIN r_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 4.000 ;
    END
  END r_data[27]
  PIN r_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END r_data[28]
  PIN r_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1931.240 4.000 1931.840 ;
    END
  END r_data[29]
  PIN r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 1996.000 1871.190 2000.000 ;
    END
  END r_data[2]
  PIN r_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END r_data[30]
  PIN r_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 425.040 2000.000 425.640 ;
    END
  END r_data[31]
  PIN r_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END r_data[32]
  PIN r_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END r_data[33]
  PIN r_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 1996.000 615.390 2000.000 ;
    END
  END r_data[34]
  PIN r_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.230 0.000 1568.510 4.000 ;
    END
  END r_data[35]
  PIN r_data[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END r_data[36]
  PIN r_data[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END r_data[37]
  PIN r_data[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 258.440 2000.000 259.040 ;
    END
  END r_data[38]
  PIN r_data[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1530.040 2000.000 1530.640 ;
    END
  END r_data[39]
  PIN r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1033.640 2000.000 1034.240 ;
    END
  END r_data[3]
  PIN r_data[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END r_data[40]
  PIN r_data[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1159.440 4.000 1160.040 ;
    END
  END r_data[41]
  PIN r_data[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 537.240 2000.000 537.840 ;
    END
  END r_data[42]
  PIN r_data[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END r_data[43]
  PIN r_data[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1200.240 2000.000 1200.840 ;
    END
  END r_data[44]
  PIN r_data[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1751.040 2000.000 1751.640 ;
    END
  END r_data[45]
  PIN r_data[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END r_data[46]
  PIN r_data[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1863.240 2000.000 1863.840 ;
    END
  END r_data[47]
  PIN r_data[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END r_data[48]
  PIN r_data[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1655.840 4.000 1656.440 ;
    END
  END r_data[49]
  PIN r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END r_data[4]
  PIN r_data[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END r_data[50]
  PIN r_data[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END r_data[51]
  PIN r_data[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END r_data[52]
  PIN r_data[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 1996.000 457.610 2000.000 ;
    END
  END r_data[53]
  PIN r_data[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 1996.000 1191.770 2000.000 ;
    END
  END r_data[54]
  PIN r_data[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.840 4.000 1435.440 ;
    END
  END r_data[55]
  PIN r_data[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END r_data[56]
  PIN r_data[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END r_data[57]
  PIN r_data[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END r_data[58]
  PIN r_data[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.230 1996.000 1085.510 2000.000 ;
    END
  END r_data[59]
  PIN r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 4.000 ;
    END
  END r_data[5]
  PIN r_data[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.650 1996.000 1764.930 2000.000 ;
    END
  END r_data[60]
  PIN r_data[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 316.240 2000.000 316.840 ;
    END
  END r_data[61]
  PIN r_data[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1822.440 4.000 1823.040 ;
    END
  END r_data[62]
  PIN r_data[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END r_data[63]
  PIN r_data[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END r_data[64]
  PIN r_data[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END r_data[65]
  PIN r_data[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END r_data[66]
  PIN r_data[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 1309.040 2000.000 1309.640 ;
    END
  END r_data[67]
  PIN r_data[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END r_data[68]
  PIN r_data[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 1996.000 1504.110 2000.000 ;
    END
  END r_data[69]
  PIN r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 1996.000 1452.590 2000.000 ;
    END
  END r_data[6]
  PIN r_data[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1996.000 39.010 2000.000 ;
    END
  END r_data[70]
  PIN r_data[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 1996.000 351.350 2000.000 ;
    END
  END r_data[71]
  PIN r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.930 0.000 1359.210 4.000 ;
    END
  END r_data[7]
  PIN r_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END r_data[8]
  PIN r_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END r_data[9]
  PIN wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 924.840 2000.000 925.440 ;
    END
  END wr
  OBS
      LAYER li1 ;
        RECT 400.200 402.475 1599.880 1599.445 ;
      LAYER met1 ;
        RECT 0.070 17.040 1987.130 1978.420 ;
      LAYER met2 ;
        RECT 0.100 1995.720 38.450 1996.210 ;
        RECT 39.290 1995.720 89.970 1996.210 ;
        RECT 90.810 1995.720 141.490 1996.210 ;
        RECT 142.330 1995.720 196.230 1996.210 ;
        RECT 197.070 1995.720 247.750 1996.210 ;
        RECT 248.590 1995.720 299.270 1996.210 ;
        RECT 300.110 1995.720 350.790 1996.210 ;
        RECT 351.630 1995.720 405.530 1996.210 ;
        RECT 406.370 1995.720 457.050 1996.210 ;
        RECT 457.890 1995.720 508.570 1996.210 ;
        RECT 509.410 1995.720 560.090 1996.210 ;
        RECT 560.930 1995.720 614.830 1996.210 ;
        RECT 615.670 1995.720 666.350 1996.210 ;
        RECT 667.190 1995.720 717.870 1996.210 ;
        RECT 718.710 1995.720 772.610 1996.210 ;
        RECT 773.450 1995.720 824.130 1996.210 ;
        RECT 824.970 1995.720 875.650 1996.210 ;
        RECT 876.490 1995.720 927.170 1996.210 ;
        RECT 928.010 1995.720 981.910 1996.210 ;
        RECT 982.750 1995.720 1033.430 1996.210 ;
        RECT 1034.270 1995.720 1084.950 1996.210 ;
        RECT 1085.790 1995.720 1136.470 1996.210 ;
        RECT 1137.310 1995.720 1191.210 1996.210 ;
        RECT 1192.050 1995.720 1242.730 1996.210 ;
        RECT 1243.570 1995.720 1294.250 1996.210 ;
        RECT 1295.090 1995.720 1345.770 1996.210 ;
        RECT 1346.610 1995.720 1400.510 1996.210 ;
        RECT 1401.350 1995.720 1452.030 1996.210 ;
        RECT 1452.870 1995.720 1503.550 1996.210 ;
        RECT 1504.390 1995.720 1555.070 1996.210 ;
        RECT 1555.910 1995.720 1609.810 1996.210 ;
        RECT 1610.650 1995.720 1661.330 1996.210 ;
        RECT 1662.170 1995.720 1712.850 1996.210 ;
        RECT 1713.690 1995.720 1764.370 1996.210 ;
        RECT 1765.210 1995.720 1819.110 1996.210 ;
        RECT 1819.950 1995.720 1870.630 1996.210 ;
        RECT 1871.470 1995.720 1922.150 1996.210 ;
        RECT 1922.990 1995.720 1973.670 1996.210 ;
        RECT 1974.510 1995.720 1987.100 1996.210 ;
        RECT 0.100 4.280 1987.100 1995.720 ;
        RECT 0.650 4.000 51.330 4.280 ;
        RECT 52.170 4.000 102.850 4.280 ;
        RECT 103.690 4.000 154.370 4.280 ;
        RECT 155.210 4.000 209.110 4.280 ;
        RECT 209.950 4.000 260.630 4.280 ;
        RECT 261.470 4.000 312.150 4.280 ;
        RECT 312.990 4.000 363.670 4.280 ;
        RECT 364.510 4.000 418.410 4.280 ;
        RECT 419.250 4.000 469.930 4.280 ;
        RECT 470.770 4.000 521.450 4.280 ;
        RECT 522.290 4.000 572.970 4.280 ;
        RECT 573.810 4.000 627.710 4.280 ;
        RECT 628.550 4.000 679.230 4.280 ;
        RECT 680.070 4.000 730.750 4.280 ;
        RECT 731.590 4.000 782.270 4.280 ;
        RECT 783.110 4.000 837.010 4.280 ;
        RECT 837.850 4.000 888.530 4.280 ;
        RECT 889.370 4.000 940.050 4.280 ;
        RECT 940.890 4.000 991.570 4.280 ;
        RECT 992.410 4.000 1046.310 4.280 ;
        RECT 1047.150 4.000 1097.830 4.280 ;
        RECT 1098.670 4.000 1149.350 4.280 ;
        RECT 1150.190 4.000 1200.870 4.280 ;
        RECT 1201.710 4.000 1255.610 4.280 ;
        RECT 1256.450 4.000 1307.130 4.280 ;
        RECT 1307.970 4.000 1358.650 4.280 ;
        RECT 1359.490 4.000 1410.170 4.280 ;
        RECT 1411.010 4.000 1464.910 4.280 ;
        RECT 1465.750 4.000 1516.430 4.280 ;
        RECT 1517.270 4.000 1567.950 4.280 ;
        RECT 1568.790 4.000 1619.470 4.280 ;
        RECT 1620.310 4.000 1674.210 4.280 ;
        RECT 1675.050 4.000 1725.730 4.280 ;
        RECT 1726.570 4.000 1777.250 4.280 ;
        RECT 1778.090 4.000 1828.770 4.280 ;
        RECT 1829.610 4.000 1883.510 4.280 ;
        RECT 1884.350 4.000 1935.030 4.280 ;
        RECT 1935.870 4.000 1986.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 1930.840 1996.000 1931.705 ;
        RECT 4.000 1918.640 1996.000 1930.840 ;
        RECT 4.000 1917.240 1995.600 1918.640 ;
        RECT 4.000 1877.840 1996.000 1917.240 ;
        RECT 4.400 1876.440 1996.000 1877.840 ;
        RECT 4.000 1864.240 1996.000 1876.440 ;
        RECT 4.000 1862.840 1995.600 1864.240 ;
        RECT 4.000 1823.440 1996.000 1862.840 ;
        RECT 4.400 1822.040 1996.000 1823.440 ;
        RECT 4.000 1809.840 1996.000 1822.040 ;
        RECT 4.000 1808.440 1995.600 1809.840 ;
        RECT 4.000 1769.040 1996.000 1808.440 ;
        RECT 4.400 1767.640 1996.000 1769.040 ;
        RECT 4.000 1752.040 1996.000 1767.640 ;
        RECT 4.000 1750.640 1995.600 1752.040 ;
        RECT 4.000 1711.240 1996.000 1750.640 ;
        RECT 4.400 1709.840 1996.000 1711.240 ;
        RECT 4.000 1697.640 1996.000 1709.840 ;
        RECT 4.000 1696.240 1995.600 1697.640 ;
        RECT 4.000 1656.840 1996.000 1696.240 ;
        RECT 4.400 1655.440 1996.000 1656.840 ;
        RECT 4.000 1643.240 1996.000 1655.440 ;
        RECT 4.000 1641.840 1995.600 1643.240 ;
        RECT 4.000 1602.440 1996.000 1641.840 ;
        RECT 4.400 1601.040 1996.000 1602.440 ;
        RECT 4.000 1588.840 1996.000 1601.040 ;
        RECT 4.000 1587.440 1995.600 1588.840 ;
        RECT 4.000 1548.040 1996.000 1587.440 ;
        RECT 4.400 1546.640 1996.000 1548.040 ;
        RECT 4.000 1531.040 1996.000 1546.640 ;
        RECT 4.000 1529.640 1995.600 1531.040 ;
        RECT 4.000 1490.240 1996.000 1529.640 ;
        RECT 4.400 1488.840 1996.000 1490.240 ;
        RECT 4.000 1476.640 1996.000 1488.840 ;
        RECT 4.000 1475.240 1995.600 1476.640 ;
        RECT 4.000 1435.840 1996.000 1475.240 ;
        RECT 4.400 1434.440 1996.000 1435.840 ;
        RECT 4.000 1422.240 1996.000 1434.440 ;
        RECT 4.000 1420.840 1995.600 1422.240 ;
        RECT 4.000 1381.440 1996.000 1420.840 ;
        RECT 4.400 1380.040 1996.000 1381.440 ;
        RECT 4.000 1367.840 1996.000 1380.040 ;
        RECT 4.000 1366.440 1995.600 1367.840 ;
        RECT 4.000 1327.040 1996.000 1366.440 ;
        RECT 4.400 1325.640 1996.000 1327.040 ;
        RECT 4.000 1310.040 1996.000 1325.640 ;
        RECT 4.000 1308.640 1995.600 1310.040 ;
        RECT 4.000 1269.240 1996.000 1308.640 ;
        RECT 4.400 1267.840 1996.000 1269.240 ;
        RECT 4.000 1255.640 1996.000 1267.840 ;
        RECT 4.000 1254.240 1995.600 1255.640 ;
        RECT 4.000 1214.840 1996.000 1254.240 ;
        RECT 4.400 1213.440 1996.000 1214.840 ;
        RECT 4.000 1201.240 1996.000 1213.440 ;
        RECT 4.000 1199.840 1995.600 1201.240 ;
        RECT 4.000 1160.440 1996.000 1199.840 ;
        RECT 4.400 1159.040 1996.000 1160.440 ;
        RECT 4.000 1146.840 1996.000 1159.040 ;
        RECT 4.000 1145.440 1995.600 1146.840 ;
        RECT 4.000 1106.040 1996.000 1145.440 ;
        RECT 4.400 1104.640 1996.000 1106.040 ;
        RECT 4.000 1089.040 1996.000 1104.640 ;
        RECT 4.000 1087.640 1995.600 1089.040 ;
        RECT 4.000 1048.240 1996.000 1087.640 ;
        RECT 4.400 1046.840 1996.000 1048.240 ;
        RECT 4.000 1034.640 1996.000 1046.840 ;
        RECT 4.000 1033.240 1995.600 1034.640 ;
        RECT 4.000 993.840 1996.000 1033.240 ;
        RECT 4.400 992.440 1996.000 993.840 ;
        RECT 4.000 980.240 1996.000 992.440 ;
        RECT 4.000 978.840 1995.600 980.240 ;
        RECT 4.000 939.440 1996.000 978.840 ;
        RECT 4.400 938.040 1996.000 939.440 ;
        RECT 4.000 925.840 1996.000 938.040 ;
        RECT 4.000 924.440 1995.600 925.840 ;
        RECT 4.000 885.040 1996.000 924.440 ;
        RECT 4.400 883.640 1996.000 885.040 ;
        RECT 4.000 868.040 1996.000 883.640 ;
        RECT 4.000 866.640 1995.600 868.040 ;
        RECT 4.000 827.240 1996.000 866.640 ;
        RECT 4.400 825.840 1996.000 827.240 ;
        RECT 4.000 813.640 1996.000 825.840 ;
        RECT 4.000 812.240 1995.600 813.640 ;
        RECT 4.000 772.840 1996.000 812.240 ;
        RECT 4.400 771.440 1996.000 772.840 ;
        RECT 4.000 759.240 1996.000 771.440 ;
        RECT 4.000 757.840 1995.600 759.240 ;
        RECT 4.000 718.440 1996.000 757.840 ;
        RECT 4.400 717.040 1996.000 718.440 ;
        RECT 4.000 704.840 1996.000 717.040 ;
        RECT 4.000 703.440 1995.600 704.840 ;
        RECT 4.000 664.040 1996.000 703.440 ;
        RECT 4.400 662.640 1996.000 664.040 ;
        RECT 4.000 647.040 1996.000 662.640 ;
        RECT 4.000 645.640 1995.600 647.040 ;
        RECT 4.000 606.240 1996.000 645.640 ;
        RECT 4.400 604.840 1996.000 606.240 ;
        RECT 4.000 592.640 1996.000 604.840 ;
        RECT 4.000 591.240 1995.600 592.640 ;
        RECT 4.000 551.840 1996.000 591.240 ;
        RECT 4.400 550.440 1996.000 551.840 ;
        RECT 4.000 538.240 1996.000 550.440 ;
        RECT 4.000 536.840 1995.600 538.240 ;
        RECT 4.000 497.440 1996.000 536.840 ;
        RECT 4.400 496.040 1996.000 497.440 ;
        RECT 4.000 480.440 1996.000 496.040 ;
        RECT 4.000 479.040 1995.600 480.440 ;
        RECT 4.000 443.040 1996.000 479.040 ;
        RECT 4.400 441.640 1996.000 443.040 ;
        RECT 4.000 426.040 1996.000 441.640 ;
        RECT 4.000 424.640 1995.600 426.040 ;
        RECT 4.000 385.240 1996.000 424.640 ;
        RECT 4.400 383.840 1996.000 385.240 ;
        RECT 4.000 371.640 1996.000 383.840 ;
        RECT 4.000 370.240 1995.600 371.640 ;
        RECT 4.000 330.840 1996.000 370.240 ;
        RECT 4.400 329.440 1996.000 330.840 ;
        RECT 4.000 317.240 1996.000 329.440 ;
        RECT 4.000 315.840 1995.600 317.240 ;
        RECT 4.000 276.440 1996.000 315.840 ;
        RECT 4.400 275.040 1996.000 276.440 ;
        RECT 4.000 259.440 1996.000 275.040 ;
        RECT 4.000 258.040 1995.600 259.440 ;
        RECT 4.000 222.040 1996.000 258.040 ;
        RECT 4.400 220.640 1996.000 222.040 ;
        RECT 4.000 205.040 1996.000 220.640 ;
        RECT 4.000 203.640 1995.600 205.040 ;
        RECT 4.000 164.240 1996.000 203.640 ;
        RECT 4.400 162.840 1996.000 164.240 ;
        RECT 4.000 150.640 1996.000 162.840 ;
        RECT 4.000 149.240 1995.600 150.640 ;
        RECT 4.000 109.840 1996.000 149.240 ;
        RECT 4.400 108.440 1996.000 109.840 ;
        RECT 4.000 96.240 1996.000 108.440 ;
        RECT 4.000 94.840 1995.600 96.240 ;
        RECT 4.000 55.440 1996.000 94.840 ;
        RECT 4.400 54.575 1996.000 55.440 ;
  END
END dff_ram
END LIBRARY

