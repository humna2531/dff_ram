magic
tech sky130A
magscale 1 2
timestamp 1709554452
<< obsli1 >>
rect 80040 80495 319976 319889
<< obsm1 >>
rect 14 3408 397426 395684
<< metal2 >>
rect 7746 399200 7802 400000
rect 18050 399200 18106 400000
rect 28354 399200 28410 400000
rect 39302 399200 39358 400000
rect 49606 399200 49662 400000
rect 59910 399200 59966 400000
rect 70214 399200 70270 400000
rect 81162 399200 81218 400000
rect 91466 399200 91522 400000
rect 101770 399200 101826 400000
rect 112074 399200 112130 400000
rect 123022 399200 123078 400000
rect 133326 399200 133382 400000
rect 143630 399200 143686 400000
rect 154578 399200 154634 400000
rect 164882 399200 164938 400000
rect 175186 399200 175242 400000
rect 185490 399200 185546 400000
rect 196438 399200 196494 400000
rect 206742 399200 206798 400000
rect 217046 399200 217102 400000
rect 227350 399200 227406 400000
rect 238298 399200 238354 400000
rect 248602 399200 248658 400000
rect 258906 399200 258962 400000
rect 269210 399200 269266 400000
rect 280158 399200 280214 400000
rect 290462 399200 290518 400000
rect 300766 399200 300822 400000
rect 311070 399200 311126 400000
rect 322018 399200 322074 400000
rect 332322 399200 332378 400000
rect 342626 399200 342682 400000
rect 352930 399200 352986 400000
rect 363878 399200 363934 400000
rect 374182 399200 374238 400000
rect 384486 399200 384542 400000
rect 394790 399200 394846 400000
rect 18 0 74 800
rect 10322 0 10378 800
rect 20626 0 20682 800
rect 30930 0 30986 800
rect 41878 0 41934 800
rect 52182 0 52238 800
rect 62486 0 62542 800
rect 72790 0 72846 800
rect 83738 0 83794 800
rect 94042 0 94098 800
rect 104346 0 104402 800
rect 114650 0 114706 800
rect 125598 0 125654 800
rect 135902 0 135958 800
rect 146206 0 146262 800
rect 156510 0 156566 800
rect 167458 0 167514 800
rect 177762 0 177818 800
rect 188066 0 188122 800
rect 198370 0 198426 800
rect 209318 0 209374 800
rect 219622 0 219678 800
rect 229926 0 229982 800
rect 240230 0 240286 800
rect 251178 0 251234 800
rect 261482 0 261538 800
rect 271786 0 271842 800
rect 282090 0 282146 800
rect 293038 0 293094 800
rect 303342 0 303398 800
rect 313646 0 313702 800
rect 323950 0 324006 800
rect 334898 0 334954 800
rect 345202 0 345258 800
rect 355506 0 355562 800
rect 365810 0 365866 800
rect 376758 0 376814 800
rect 387062 0 387118 800
rect 397366 0 397422 800
<< obsm2 >>
rect 20 399144 7690 399242
rect 7858 399144 17994 399242
rect 18162 399144 28298 399242
rect 28466 399144 39246 399242
rect 39414 399144 49550 399242
rect 49718 399144 59854 399242
rect 60022 399144 70158 399242
rect 70326 399144 81106 399242
rect 81274 399144 91410 399242
rect 91578 399144 101714 399242
rect 101882 399144 112018 399242
rect 112186 399144 122966 399242
rect 123134 399144 133270 399242
rect 133438 399144 143574 399242
rect 143742 399144 154522 399242
rect 154690 399144 164826 399242
rect 164994 399144 175130 399242
rect 175298 399144 185434 399242
rect 185602 399144 196382 399242
rect 196550 399144 206686 399242
rect 206854 399144 216990 399242
rect 217158 399144 227294 399242
rect 227462 399144 238242 399242
rect 238410 399144 248546 399242
rect 248714 399144 258850 399242
rect 259018 399144 269154 399242
rect 269322 399144 280102 399242
rect 280270 399144 290406 399242
rect 290574 399144 300710 399242
rect 300878 399144 311014 399242
rect 311182 399144 321962 399242
rect 322130 399144 332266 399242
rect 332434 399144 342570 399242
rect 342738 399144 352874 399242
rect 353042 399144 363822 399242
rect 363990 399144 374126 399242
rect 374294 399144 384430 399242
rect 384598 399144 394734 399242
rect 394902 399144 397420 399242
rect 20 856 397420 399144
rect 130 800 10266 856
rect 10434 800 20570 856
rect 20738 800 30874 856
rect 31042 800 41822 856
rect 41990 800 52126 856
rect 52294 800 62430 856
rect 62598 800 72734 856
rect 72902 800 83682 856
rect 83850 800 93986 856
rect 94154 800 104290 856
rect 104458 800 114594 856
rect 114762 800 125542 856
rect 125710 800 135846 856
rect 136014 800 146150 856
rect 146318 800 156454 856
rect 156622 800 167402 856
rect 167570 800 177706 856
rect 177874 800 188010 856
rect 188178 800 198314 856
rect 198482 800 209262 856
rect 209430 800 219566 856
rect 219734 800 229870 856
rect 230038 800 240174 856
rect 240342 800 251122 856
rect 251290 800 261426 856
rect 261594 800 271730 856
rect 271898 800 282034 856
rect 282202 800 292982 856
rect 293150 800 303286 856
rect 303454 800 313590 856
rect 313758 800 323894 856
rect 324062 800 334842 856
rect 335010 800 345146 856
rect 345314 800 355450 856
rect 355618 800 365754 856
rect 365922 800 376702 856
rect 376870 800 387006 856
rect 387174 800 397310 856
<< metal3 >>
rect 0 397808 800 397928
rect 399200 394408 400000 394528
rect 0 386248 800 386368
rect 399200 383528 400000 383648
rect 0 375368 800 375488
rect 399200 372648 400000 372768
rect 0 364488 800 364608
rect 399200 361768 400000 361888
rect 0 353608 800 353728
rect 399200 350208 400000 350328
rect 0 342048 800 342168
rect 399200 339328 400000 339448
rect 0 331168 800 331288
rect 399200 328448 400000 328568
rect 0 320288 800 320408
rect 399200 317568 400000 317688
rect 0 309408 800 309528
rect 399200 306008 400000 306128
rect 0 297848 800 297968
rect 399200 295128 400000 295248
rect 0 286968 800 287088
rect 399200 284248 400000 284368
rect 0 276088 800 276208
rect 399200 273368 400000 273488
rect 0 265208 800 265328
rect 399200 261808 400000 261928
rect 0 253648 800 253768
rect 399200 250928 400000 251048
rect 0 242768 800 242888
rect 399200 240048 400000 240168
rect 0 231888 800 232008
rect 399200 229168 400000 229288
rect 0 221008 800 221128
rect 399200 217608 400000 217728
rect 0 209448 800 209568
rect 399200 206728 400000 206848
rect 0 198568 800 198688
rect 399200 195848 400000 195968
rect 0 187688 800 187808
rect 399200 184968 400000 185088
rect 0 176808 800 176928
rect 399200 173408 400000 173528
rect 0 165248 800 165368
rect 399200 162528 400000 162648
rect 0 154368 800 154488
rect 399200 151648 400000 151768
rect 0 143488 800 143608
rect 399200 140768 400000 140888
rect 0 132608 800 132728
rect 399200 129208 400000 129328
rect 0 121048 800 121168
rect 399200 118328 400000 118448
rect 0 110168 800 110288
rect 399200 107448 400000 107568
rect 0 99288 800 99408
rect 399200 95888 400000 96008
rect 0 88408 800 88528
rect 399200 85008 400000 85128
rect 0 76848 800 76968
rect 399200 74128 400000 74248
rect 0 65968 800 66088
rect 399200 63248 400000 63368
rect 0 55088 800 55208
rect 399200 51688 400000 51808
rect 0 44208 800 44328
rect 399200 40808 400000 40928
rect 0 32648 800 32768
rect 399200 29928 400000 30048
rect 0 21768 800 21888
rect 399200 19048 400000 19168
rect 0 10888 800 11008
rect 399200 7488 400000 7608
<< obsm3 >>
rect 880 386168 399200 386341
rect 800 383728 399200 386168
rect 800 383448 399120 383728
rect 800 375568 399200 383448
rect 880 375288 399200 375568
rect 800 372848 399200 375288
rect 800 372568 399120 372848
rect 800 364688 399200 372568
rect 880 364408 399200 364688
rect 800 361968 399200 364408
rect 800 361688 399120 361968
rect 800 353808 399200 361688
rect 880 353528 399200 353808
rect 800 350408 399200 353528
rect 800 350128 399120 350408
rect 800 342248 399200 350128
rect 880 341968 399200 342248
rect 800 339528 399200 341968
rect 800 339248 399120 339528
rect 800 331368 399200 339248
rect 880 331088 399200 331368
rect 800 328648 399200 331088
rect 800 328368 399120 328648
rect 800 320488 399200 328368
rect 880 320208 399200 320488
rect 800 317768 399200 320208
rect 800 317488 399120 317768
rect 800 309608 399200 317488
rect 880 309328 399200 309608
rect 800 306208 399200 309328
rect 800 305928 399120 306208
rect 800 298048 399200 305928
rect 880 297768 399200 298048
rect 800 295328 399200 297768
rect 800 295048 399120 295328
rect 800 287168 399200 295048
rect 880 286888 399200 287168
rect 800 284448 399200 286888
rect 800 284168 399120 284448
rect 800 276288 399200 284168
rect 880 276008 399200 276288
rect 800 273568 399200 276008
rect 800 273288 399120 273568
rect 800 265408 399200 273288
rect 880 265128 399200 265408
rect 800 262008 399200 265128
rect 800 261728 399120 262008
rect 800 253848 399200 261728
rect 880 253568 399200 253848
rect 800 251128 399200 253568
rect 800 250848 399120 251128
rect 800 242968 399200 250848
rect 880 242688 399200 242968
rect 800 240248 399200 242688
rect 800 239968 399120 240248
rect 800 232088 399200 239968
rect 880 231808 399200 232088
rect 800 229368 399200 231808
rect 800 229088 399120 229368
rect 800 221208 399200 229088
rect 880 220928 399200 221208
rect 800 217808 399200 220928
rect 800 217528 399120 217808
rect 800 209648 399200 217528
rect 880 209368 399200 209648
rect 800 206928 399200 209368
rect 800 206648 399120 206928
rect 800 198768 399200 206648
rect 880 198488 399200 198768
rect 800 196048 399200 198488
rect 800 195768 399120 196048
rect 800 187888 399200 195768
rect 880 187608 399200 187888
rect 800 185168 399200 187608
rect 800 184888 399120 185168
rect 800 177008 399200 184888
rect 880 176728 399200 177008
rect 800 173608 399200 176728
rect 800 173328 399120 173608
rect 800 165448 399200 173328
rect 880 165168 399200 165448
rect 800 162728 399200 165168
rect 800 162448 399120 162728
rect 800 154568 399200 162448
rect 880 154288 399200 154568
rect 800 151848 399200 154288
rect 800 151568 399120 151848
rect 800 143688 399200 151568
rect 880 143408 399200 143688
rect 800 140968 399200 143408
rect 800 140688 399120 140968
rect 800 132808 399200 140688
rect 880 132528 399200 132808
rect 800 129408 399200 132528
rect 800 129128 399120 129408
rect 800 121248 399200 129128
rect 880 120968 399200 121248
rect 800 118528 399200 120968
rect 800 118248 399120 118528
rect 800 110368 399200 118248
rect 880 110088 399200 110368
rect 800 107648 399200 110088
rect 800 107368 399120 107648
rect 800 99488 399200 107368
rect 880 99208 399200 99488
rect 800 96088 399200 99208
rect 800 95808 399120 96088
rect 800 88608 399200 95808
rect 880 88328 399200 88608
rect 800 85208 399200 88328
rect 800 84928 399120 85208
rect 800 77048 399200 84928
rect 880 76768 399200 77048
rect 800 74328 399200 76768
rect 800 74048 399120 74328
rect 800 66168 399200 74048
rect 880 65888 399200 66168
rect 800 63448 399200 65888
rect 800 63168 399120 63448
rect 800 55288 399200 63168
rect 880 55008 399200 55288
rect 800 51888 399200 55008
rect 800 51608 399120 51888
rect 800 44408 399200 51608
rect 880 44128 399200 44408
rect 800 41008 399200 44128
rect 800 40728 399120 41008
rect 800 32848 399200 40728
rect 880 32568 399200 32848
rect 800 30128 399200 32568
rect 800 29848 399120 30128
rect 800 21968 399200 29848
rect 880 21688 399200 21968
rect 800 19248 399200 21688
rect 800 18968 399120 19248
rect 800 11088 399200 18968
rect 880 10915 399200 11088
<< metal4 >>
rect 83144 80464 83464 319920
rect 83804 80464 84124 319920
rect 113864 80464 114184 319920
rect 114524 80464 114844 319920
rect 144584 80464 144904 319920
rect 145244 80464 145564 319920
rect 175304 80464 175624 319920
rect 175964 80464 176284 319920
rect 206024 80464 206344 319920
rect 206684 80464 207004 319920
rect 236744 80464 237064 319920
rect 237404 80464 237724 319920
rect 267464 80464 267784 319920
rect 268124 80464 268444 319920
rect 298184 80464 298504 319920
rect 298844 80464 299164 319920
<< metal5 >>
rect 79992 298794 320024 299114
rect 79992 298134 320024 298454
rect 79992 268158 320024 268478
rect 79992 267498 320024 267818
rect 79992 237522 320024 237842
rect 79992 236862 320024 237182
rect 79992 206886 320024 207206
rect 79992 206226 320024 206546
rect 79992 176250 320024 176570
rect 79992 175590 320024 175910
rect 79992 145614 320024 145934
rect 79992 144954 320024 145274
rect 79992 114978 320024 115298
rect 79992 114318 320024 114638
rect 79992 84342 320024 84662
rect 79992 83682 320024 84002
<< labels >>
rlabel metal4 s 83804 80464 84124 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 114524 80464 114844 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 145244 80464 145564 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 175964 80464 176284 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 206684 80464 207004 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 237404 80464 237724 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 268124 80464 268444 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298844 80464 299164 319920 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 84342 320024 84662 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 114978 320024 115298 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 145614 320024 145934 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 176250 320024 176570 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 206886 320024 207206 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 237522 320024 237842 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 268158 320024 268478 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 79992 298794 320024 299114 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 83144 80464 83464 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 113864 80464 114184 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 144584 80464 144904 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 175304 80464 175624 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 206024 80464 206344 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 236744 80464 237064 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 267464 80464 267784 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 298184 80464 298504 319920 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 83682 320024 84002 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 114318 320024 114638 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 144954 320024 145274 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 175590 320024 175910 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 206226 320024 206546 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 236862 320024 237182 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 267498 320024 267818 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 79992 298134 320024 298454 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 196438 399200 196494 400000 6 addr[0]
port 3 nsew signal input
rlabel metal3 s 0 297848 800 297968 6 addr[1]
port 4 nsew signal input
rlabel metal3 s 0 132608 800 132728 6 clk
port 5 nsew signal input
rlabel metal3 s 399200 129208 400000 129328 6 data[0]
port 6 nsew signal input
rlabel metal3 s 399200 151648 400000 151768 6 data[10]
port 7 nsew signal input
rlabel metal3 s 0 320288 800 320408 6 data[11]
port 8 nsew signal input
rlabel metal2 s 28354 399200 28410 400000 6 data[12]
port 9 nsew signal input
rlabel metal2 s 133326 399200 133382 400000 6 data[13]
port 10 nsew signal input
rlabel metal2 s 355506 0 355562 800 6 data[14]
port 11 nsew signal input
rlabel metal2 s 164882 399200 164938 400000 6 data[15]
port 12 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 data[16]
port 13 nsew signal input
rlabel metal2 s 206742 399200 206798 400000 6 data[17]
port 14 nsew signal input
rlabel metal3 s 0 397808 800 397928 6 data[18]
port 15 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 data[19]
port 16 nsew signal input
rlabel metal2 s 175186 399200 175242 400000 6 data[1]
port 17 nsew signal input
rlabel metal2 s 49606 399200 49662 400000 6 data[20]
port 18 nsew signal input
rlabel metal3 s 399200 284248 400000 284368 6 data[21]
port 19 nsew signal input
rlabel metal3 s 0 265208 800 265328 6 data[22]
port 20 nsew signal input
rlabel metal3 s 0 375368 800 375488 6 data[23]
port 21 nsew signal input
rlabel metal2 s 112074 399200 112130 400000 6 data[24]
port 22 nsew signal input
rlabel metal3 s 0 221008 800 221128 6 data[25]
port 23 nsew signal input
rlabel metal3 s 0 342048 800 342168 6 data[26]
port 24 nsew signal input
rlabel metal3 s 399200 328448 400000 328568 6 data[27]
port 25 nsew signal input
rlabel metal3 s 399200 217608 400000 217728 6 data[28]
port 26 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 data[29]
port 27 nsew signal input
rlabel metal2 s 280158 399200 280214 400000 6 data[2]
port 28 nsew signal input
rlabel metal3 s 399200 394408 400000 394528 6 data[30]
port 29 nsew signal input
rlabel metal3 s 399200 317568 400000 317688 6 data[31]
port 30 nsew signal input
rlabel metal3 s 399200 162528 400000 162648 6 data[32]
port 31 nsew signal input
rlabel metal2 s 261482 0 261538 800 6 data[33]
port 32 nsew signal input
rlabel metal2 s 269210 399200 269266 400000 6 data[34]
port 33 nsew signal input
rlabel metal2 s 332322 399200 332378 400000 6 data[35]
port 34 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 data[36]
port 35 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 data[37]
port 36 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 data[38]
port 37 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 data[39]
port 38 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 data[3]
port 39 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 data[40]
port 40 nsew signal input
rlabel metal3 s 0 253648 800 253768 6 data[41]
port 41 nsew signal input
rlabel metal3 s 399200 140768 400000 140888 6 data[42]
port 42 nsew signal input
rlabel metal3 s 399200 250928 400000 251048 6 data[43]
port 43 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 data[44]
port 44 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 data[45]
port 45 nsew signal input
rlabel metal3 s 399200 195848 400000 195968 6 data[46]
port 46 nsew signal input
rlabel metal2 s 227350 399200 227406 400000 6 data[47]
port 47 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 data[48]
port 48 nsew signal input
rlabel metal2 s 185490 399200 185546 400000 6 data[49]
port 49 nsew signal input
rlabel metal3 s 399200 19048 400000 19168 6 data[4]
port 50 nsew signal input
rlabel metal3 s 399200 339328 400000 339448 6 data[50]
port 51 nsew signal input
rlabel metal2 s 394790 399200 394846 400000 6 data[51]
port 52 nsew signal input
rlabel metal2 s 143630 399200 143686 400000 6 data[52]
port 53 nsew signal input
rlabel metal2 s 303342 0 303398 800 6 data[53]
port 54 nsew signal input
rlabel metal3 s 399200 295128 400000 295248 6 data[54]
port 55 nsew signal input
rlabel metal2 s 342626 399200 342682 400000 6 data[55]
port 56 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 data[56]
port 57 nsew signal input
rlabel metal2 s 384486 399200 384542 400000 6 data[57]
port 58 nsew signal input
rlabel metal3 s 399200 361768 400000 361888 6 data[58]
port 59 nsew signal input
rlabel metal2 s 59910 399200 59966 400000 6 data[59]
port 60 nsew signal input
rlabel metal3 s 399200 7488 400000 7608 6 data[5]
port 61 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 data[60]
port 62 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 data[61]
port 63 nsew signal input
rlabel metal2 s 251178 0 251234 800 6 data[62]
port 64 nsew signal input
rlabel metal2 s 39302 399200 39358 400000 6 data[63]
port 65 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 data[64]
port 66 nsew signal input
rlabel metal2 s 18050 399200 18106 400000 6 data[65]
port 67 nsew signal input
rlabel metal2 s 258906 399200 258962 400000 6 data[66]
port 68 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 data[67]
port 69 nsew signal input
rlabel metal3 s 399200 29928 400000 30048 6 data[68]
port 70 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 data[69]
port 71 nsew signal input
rlabel metal3 s 399200 95888 400000 96008 6 data[6]
port 72 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 data[70]
port 73 nsew signal input
rlabel metal3 s 399200 383528 400000 383648 6 data[71]
port 74 nsew signal input
rlabel metal3 s 399200 118328 400000 118448 6 data[7]
port 75 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 data[8]
port 76 nsew signal input
rlabel metal3 s 0 242768 800 242888 6 data[9]
port 77 nsew signal input
rlabel metal2 s 311070 399200 311126 400000 6 enb
port 78 nsew signal input
rlabel metal2 s 101770 399200 101826 400000 6 r_data[0]
port 79 nsew signal output
rlabel metal3 s 0 276088 800 276208 6 r_data[10]
port 80 nsew signal output
rlabel metal3 s 399200 273368 400000 273488 6 r_data[11]
port 81 nsew signal output
rlabel metal3 s 399200 74128 400000 74248 6 r_data[12]
port 82 nsew signal output
rlabel metal2 s 322018 399200 322074 400000 6 r_data[13]
port 83 nsew signal output
rlabel metal2 s 248602 399200 248658 400000 6 r_data[14]
port 84 nsew signal output
rlabel metal2 s 363878 399200 363934 400000 6 r_data[15]
port 85 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 r_data[16]
port 86 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 r_data[17]
port 87 nsew signal output
rlabel metal2 s 397366 0 397422 800 6 r_data[18]
port 88 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 r_data[19]
port 89 nsew signal output
rlabel metal3 s 399200 229168 400000 229288 6 r_data[1]
port 90 nsew signal output
rlabel metal3 s 399200 173408 400000 173528 6 r_data[20]
port 91 nsew signal output
rlabel metal2 s 154578 399200 154634 400000 6 r_data[21]
port 92 nsew signal output
rlabel metal2 s 81162 399200 81218 400000 6 r_data[22]
port 93 nsew signal output
rlabel metal3 s 399200 40808 400000 40928 6 r_data[23]
port 94 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 r_data[24]
port 95 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 r_data[25]
port 96 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 r_data[26]
port 97 nsew signal output
rlabel metal2 s 376758 0 376814 800 6 r_data[27]
port 98 nsew signal output
rlabel metal2 s 198370 0 198426 800 6 r_data[28]
port 99 nsew signal output
rlabel metal3 s 0 386248 800 386368 6 r_data[29]
port 100 nsew signal output
rlabel metal2 s 374182 399200 374238 400000 6 r_data[2]
port 101 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 r_data[30]
port 102 nsew signal output
rlabel metal3 s 399200 85008 400000 85128 6 r_data[31]
port 103 nsew signal output
rlabel metal2 s 240230 0 240286 800 6 r_data[32]
port 104 nsew signal output
rlabel metal2 s 387062 0 387118 800 6 r_data[33]
port 105 nsew signal output
rlabel metal2 s 123022 399200 123078 400000 6 r_data[34]
port 106 nsew signal output
rlabel metal2 s 313646 0 313702 800 6 r_data[35]
port 107 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 r_data[36]
port 108 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 r_data[37]
port 109 nsew signal output
rlabel metal3 s 399200 51688 400000 51808 6 r_data[38]
port 110 nsew signal output
rlabel metal3 s 399200 306008 400000 306128 6 r_data[39]
port 111 nsew signal output
rlabel metal3 s 399200 206728 400000 206848 6 r_data[3]
port 112 nsew signal output
rlabel metal2 s 334898 0 334954 800 6 r_data[40]
port 113 nsew signal output
rlabel metal3 s 0 231888 800 232008 6 r_data[41]
port 114 nsew signal output
rlabel metal3 s 399200 107448 400000 107568 6 r_data[42]
port 115 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 r_data[43]
port 116 nsew signal output
rlabel metal3 s 399200 240048 400000 240168 6 r_data[44]
port 117 nsew signal output
rlabel metal3 s 399200 350208 400000 350328 6 r_data[45]
port 118 nsew signal output
rlabel metal2 s 365810 0 365866 800 6 r_data[46]
port 119 nsew signal output
rlabel metal3 s 399200 372648 400000 372768 6 r_data[47]
port 120 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 r_data[48]
port 121 nsew signal output
rlabel metal3 s 0 331168 800 331288 6 r_data[49]
port 122 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 r_data[4]
port 123 nsew signal output
rlabel metal2 s 18 0 74 800 6 r_data[50]
port 124 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 r_data[51]
port 125 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 r_data[52]
port 126 nsew signal output
rlabel metal2 s 91466 399200 91522 400000 6 r_data[53]
port 127 nsew signal output
rlabel metal2 s 238298 399200 238354 400000 6 r_data[54]
port 128 nsew signal output
rlabel metal3 s 0 286968 800 287088 6 r_data[55]
port 129 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 r_data[56]
port 130 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 r_data[57]
port 131 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 r_data[58]
port 132 nsew signal output
rlabel metal2 s 217046 399200 217102 400000 6 r_data[59]
port 133 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 r_data[5]
port 134 nsew signal output
rlabel metal2 s 352930 399200 352986 400000 6 r_data[60]
port 135 nsew signal output
rlabel metal3 s 399200 63248 400000 63368 6 r_data[61]
port 136 nsew signal output
rlabel metal3 s 0 364488 800 364608 6 r_data[62]
port 137 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 r_data[63]
port 138 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 r_data[64]
port 139 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 r_data[65]
port 140 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 r_data[66]
port 141 nsew signal output
rlabel metal3 s 399200 261808 400000 261928 6 r_data[67]
port 142 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 r_data[68]
port 143 nsew signal output
rlabel metal2 s 300766 399200 300822 400000 6 r_data[69]
port 144 nsew signal output
rlabel metal2 s 290462 399200 290518 400000 6 r_data[6]
port 145 nsew signal output
rlabel metal2 s 7746 399200 7802 400000 6 r_data[70]
port 146 nsew signal output
rlabel metal2 s 70214 399200 70270 400000 6 r_data[71]
port 147 nsew signal output
rlabel metal2 s 271786 0 271842 800 6 r_data[7]
port 148 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 r_data[8]
port 149 nsew signal output
rlabel metal3 s 0 353608 800 353728 6 r_data[9]
port 150 nsew signal output
rlabel metal3 s 399200 184968 400000 185088 6 wr
port 151 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 400000 400000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15531218
string GDS_FILE /openlane/designs/dff_ram/runs/second_run/results/signoff/dff_ram.magic.gds
string GDS_START 197634
<< end >>

