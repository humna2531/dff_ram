module dff_ram (clk,
    enb,
    wr,
    addr,
    data,
    r_data);
 input clk;
 input enb;
 input wr;
 input [1:0] addr;
 input [71:0] data;
 output [71:0] r_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net14;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net15;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net16;
 wire net80;
 wire clknet_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__and4bb_2 _049_ (.A_N(net1),
    .B_N(net2),
    .C(net7),
    .D(net8),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _050_ (.A0(\mem[0][0] ),
    .A1(net3),
    .S(_020_),
    .X(_021_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _051_ (.A(_021_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _052_ (.A0(\mem[0][1] ),
    .A1(net4),
    .S(_020_),
    .X(_022_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _053_ (.A(_022_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _054_ (.A0(\mem[0][2] ),
    .A1(net5),
    .S(_020_),
    .X(_023_));
 sky130_fd_sc_hd__clkbuf_2 _055_ (.A(_023_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _056_ (.A0(\mem[0][3] ),
    .A1(net6),
    .S(_020_),
    .X(_024_));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(_024_),
    .X(_003_));
 sky130_fd_sc_hd__and4b_4 _058_ (.A_N(net1),
    .B(net2),
    .C(net7),
    .D(net8),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _059_ (.A0(\mem[2][0] ),
    .A1(net3),
    .S(_025_),
    .X(_026_));
 sky130_fd_sc_hd__clkbuf_2 _060_ (.A(_026_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _061_ (.A0(\mem[2][1] ),
    .A1(net4),
    .S(_025_),
    .X(_027_));
 sky130_fd_sc_hd__clkbuf_1 _062_ (.A(_027_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _063_ (.A0(\mem[2][2] ),
    .A1(net5),
    .S(_025_),
    .X(_028_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _064_ (.A(_028_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _065_ (.A0(\mem[2][3] ),
    .A1(net6),
    .S(_025_),
    .X(_029_));
 sky130_fd_sc_hd__clkbuf_1 _066_ (.A(_029_),
    .X(_007_));
 sky130_fd_sc_hd__and4b_4 _067_ (.A_N(net2),
    .B(net1),
    .C(net8),
    .D(net7),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(\mem[1][0] ),
    .A1(net3),
    .S(_030_),
    .X(_031_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _069_ (.A(_031_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _070_ (.A0(\mem[1][1] ),
    .A1(net4),
    .S(_030_),
    .X(_032_));
 sky130_fd_sc_hd__clkbuf_2 _071_ (.A(_032_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _072_ (.A0(\mem[1][2] ),
    .A1(net5),
    .S(_030_),
    .X(_033_));
 sky130_fd_sc_hd__clkbuf_2 _073_ (.A(_033_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(\mem[1][3] ),
    .A1(net6),
    .S(_030_),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(_034_),
    .X(_011_));
 sky130_fd_sc_hd__mux4_2 _076_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[2][0] ),
    .A3(\mem[3][0] ),
    .S0(net1),
    .S1(net2),
    .X(_035_));
 sky130_fd_sc_hd__and2b_2 _077_ (.A_N(net8),
    .B(net7),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(net9),
    .A1(_035_),
    .S(_036_),
    .X(_037_));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(_037_),
    .X(_012_));
 sky130_fd_sc_hd__mux4_1 _080_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[2][1] ),
    .A3(\mem[3][1] ),
    .S0(net1),
    .S1(net2),
    .X(_038_));
 sky130_fd_sc_hd__mux2_2 _081_ (.A0(net10),
    .A1(_038_),
    .S(_036_),
    .X(_039_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _082_ (.A(_039_),
    .X(_013_));
 sky130_fd_sc_hd__mux4_1 _083_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[2][2] ),
    .A3(\mem[3][2] ),
    .S0(net1),
    .S1(net2),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _084_ (.A0(net11),
    .A1(_040_),
    .S(_036_),
    .X(_041_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _085_ (.A(_041_),
    .X(_014_));
 sky130_fd_sc_hd__mux4_1 _086_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[2][3] ),
    .A3(\mem[3][3] ),
    .S0(net1),
    .S1(net2),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _087_ (.A0(net12),
    .A1(_042_),
    .S(_036_),
    .X(_043_));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(_043_),
    .X(_015_));
 sky130_fd_sc_hd__and4_4 _089_ (.A(net7),
    .B(net8),
    .C(net1),
    .D(net2),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _090_ (.A0(\mem[3][0] ),
    .A1(net3),
    .S(_044_),
    .X(_045_));
 sky130_fd_sc_hd__clkbuf_2 _091_ (.A(_045_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _092_ (.A0(\mem[3][1] ),
    .A1(net4),
    .S(_044_),
    .X(_046_));
 sky130_fd_sc_hd__clkbuf_2 _093_ (.A(_046_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _094_ (.A0(\mem[3][2] ),
    .A1(net5),
    .S(_044_),
    .X(_047_));
 sky130_fd_sc_hd__clkbuf_2 _095_ (.A(_047_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _096_ (.A0(\mem[3][3] ),
    .A1(net6),
    .S(_044_),
    .X(_048_));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(_048_),
    .X(_019_));
 sky130_fd_sc_hd__dfxtp_1 _098_ (.CLK(clknet_1_1__leaf_clk),
    .D(_000_),
    .Q(\mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _099_ (.CLK(clknet_1_1__leaf_clk),
    .D(_001_),
    .Q(\mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _100_ (.CLK(clknet_1_0__leaf_clk),
    .D(_002_),
    .Q(\mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _101_ (.CLK(clknet_1_1__leaf_clk),
    .D(_003_),
    .Q(\mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _102_ (.CLK(clknet_1_1__leaf_clk),
    .D(_004_),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_2 _103_ (.CLK(clknet_1_0__leaf_clk),
    .D(_005_),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _104_ (.CLK(clknet_1_1__leaf_clk),
    .D(_006_),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _105_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _106_ (.CLK(clknet_1_1__leaf_clk),
    .D(_008_),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_2 _107_ (.CLK(clknet_1_0__leaf_clk),
    .D(_009_),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _108_ (.CLK(clknet_1_0__leaf_clk),
    .D(_010_),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _109_ (.CLK(clknet_1_0__leaf_clk),
    .D(_011_),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_4 _110_ (.CLK(clknet_1_1__leaf_clk),
    .D(_012_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_4 _111_ (.CLK(clknet_1_1__leaf_clk),
    .D(_013_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_4 _112_ (.CLK(clknet_1_0__leaf_clk),
    .D(_014_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_4 _113_ (.CLK(clknet_1_1__leaf_clk),
    .D(_015_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _114_ (.CLK(clknet_1_1__leaf_clk),
    .D(_016_),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _115_ (.CLK(clknet_1_0__leaf_clk),
    .D(_017_),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _116_ (.CLK(clknet_1_0__leaf_clk),
    .D(_018_),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_2 _117_ (.CLK(clknet_1_1__leaf_clk),
    .D(_019_),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__conb_1 dff_ram_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 dff_ram_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 dff_ram_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 dff_ram_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 dff_ram_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 dff_ram_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 dff_ram_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 dff_ram_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 dff_ram_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 dff_ram_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 dff_ram_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 dff_ram_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 dff_ram_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 dff_ram_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 dff_ram_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 dff_ram_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 dff_ram_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 dff_ram_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 dff_ram_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 dff_ram_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 dff_ram_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 dff_ram_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 dff_ram_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 dff_ram_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 dff_ram_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 dff_ram_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 dff_ram_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 dff_ram_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 dff_ram_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 dff_ram_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 dff_ram_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 dff_ram_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 dff_ram_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 dff_ram_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 dff_ram_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 dff_ram_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 dff_ram_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 dff_ram_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 dff_ram_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 dff_ram_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 dff_ram_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 dff_ram_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 dff_ram_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 dff_ram_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 dff_ram_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 dff_ram_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 dff_ram_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 dff_ram_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 dff_ram_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 dff_ram_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 dff_ram_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 dff_ram_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 dff_ram_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 dff_ram_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 dff_ram_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 dff_ram_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 dff_ram_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 dff_ram_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 dff_ram_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 dff_ram_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 dff_ram_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 dff_ram_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 dff_ram_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 dff_ram_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 dff_ram_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 dff_ram_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 dff_ram_80 (.LO(net80));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__decap_3 PHY_644 ();
 sky130_fd_sc_hd__decap_3 PHY_645 ();
 sky130_fd_sc_hd__decap_3 PHY_646 ();
 sky130_fd_sc_hd__decap_3 PHY_647 ();
 sky130_fd_sc_hd__decap_3 PHY_648 ();
 sky130_fd_sc_hd__decap_3 PHY_649 ();
 sky130_fd_sc_hd__decap_3 PHY_650 ();
 sky130_fd_sc_hd__decap_3 PHY_651 ();
 sky130_fd_sc_hd__decap_3 PHY_652 ();
 sky130_fd_sc_hd__decap_3 PHY_653 ();
 sky130_fd_sc_hd__decap_3 PHY_654 ();
 sky130_fd_sc_hd__decap_3 PHY_655 ();
 sky130_fd_sc_hd__decap_3 PHY_656 ();
 sky130_fd_sc_hd__decap_3 PHY_657 ();
 sky130_fd_sc_hd__decap_3 PHY_658 ();
 sky130_fd_sc_hd__decap_3 PHY_659 ();
 sky130_fd_sc_hd__decap_3 PHY_660 ();
 sky130_fd_sc_hd__decap_3 PHY_661 ();
 sky130_fd_sc_hd__decap_3 PHY_662 ();
 sky130_fd_sc_hd__decap_3 PHY_663 ();
 sky130_fd_sc_hd__decap_3 PHY_664 ();
 sky130_fd_sc_hd__decap_3 PHY_665 ();
 sky130_fd_sc_hd__decap_3 PHY_666 ();
 sky130_fd_sc_hd__decap_3 PHY_667 ();
 sky130_fd_sc_hd__decap_3 PHY_668 ();
 sky130_fd_sc_hd__decap_3 PHY_669 ();
 sky130_fd_sc_hd__decap_3 PHY_670 ();
 sky130_fd_sc_hd__decap_3 PHY_671 ();
 sky130_fd_sc_hd__decap_3 PHY_672 ();
 sky130_fd_sc_hd__decap_3 PHY_673 ();
 sky130_fd_sc_hd__decap_3 PHY_674 ();
 sky130_fd_sc_hd__decap_3 PHY_675 ();
 sky130_fd_sc_hd__decap_3 PHY_676 ();
 sky130_fd_sc_hd__decap_3 PHY_677 ();
 sky130_fd_sc_hd__decap_3 PHY_678 ();
 sky130_fd_sc_hd__decap_3 PHY_679 ();
 sky130_fd_sc_hd__decap_3 PHY_680 ();
 sky130_fd_sc_hd__decap_3 PHY_681 ();
 sky130_fd_sc_hd__decap_3 PHY_682 ();
 sky130_fd_sc_hd__decap_3 PHY_683 ();
 sky130_fd_sc_hd__decap_3 PHY_684 ();
 sky130_fd_sc_hd__decap_3 PHY_685 ();
 sky130_fd_sc_hd__decap_3 PHY_686 ();
 sky130_fd_sc_hd__decap_3 PHY_687 ();
 sky130_fd_sc_hd__decap_3 PHY_688 ();
 sky130_fd_sc_hd__decap_3 PHY_689 ();
 sky130_fd_sc_hd__decap_3 PHY_690 ();
 sky130_fd_sc_hd__decap_3 PHY_691 ();
 sky130_fd_sc_hd__decap_3 PHY_692 ();
 sky130_fd_sc_hd__decap_3 PHY_693 ();
 sky130_fd_sc_hd__decap_3 PHY_694 ();
 sky130_fd_sc_hd__decap_3 PHY_695 ();
 sky130_fd_sc_hd__decap_3 PHY_696 ();
 sky130_fd_sc_hd__decap_3 PHY_697 ();
 sky130_fd_sc_hd__decap_3 PHY_698 ();
 sky130_fd_sc_hd__decap_3 PHY_699 ();
 sky130_fd_sc_hd__decap_3 PHY_700 ();
 sky130_fd_sc_hd__decap_3 PHY_701 ();
 sky130_fd_sc_hd__decap_3 PHY_702 ();
 sky130_fd_sc_hd__decap_3 PHY_703 ();
 sky130_fd_sc_hd__decap_3 PHY_704 ();
 sky130_fd_sc_hd__decap_3 PHY_705 ();
 sky130_fd_sc_hd__decap_3 PHY_706 ();
 sky130_fd_sc_hd__decap_3 PHY_707 ();
 sky130_fd_sc_hd__decap_3 PHY_708 ();
 sky130_fd_sc_hd__decap_3 PHY_709 ();
 sky130_fd_sc_hd__decap_3 PHY_710 ();
 sky130_fd_sc_hd__decap_3 PHY_711 ();
 sky130_fd_sc_hd__decap_3 PHY_712 ();
 sky130_fd_sc_hd__decap_3 PHY_713 ();
 sky130_fd_sc_hd__decap_3 PHY_714 ();
 sky130_fd_sc_hd__decap_3 PHY_715 ();
 sky130_fd_sc_hd__decap_3 PHY_716 ();
 sky130_fd_sc_hd__decap_3 PHY_717 ();
 sky130_fd_sc_hd__decap_3 PHY_718 ();
 sky130_fd_sc_hd__decap_3 PHY_719 ();
 sky130_fd_sc_hd__decap_3 PHY_720 ();
 sky130_fd_sc_hd__decap_3 PHY_721 ();
 sky130_fd_sc_hd__decap_3 PHY_722 ();
 sky130_fd_sc_hd__decap_3 PHY_723 ();
 sky130_fd_sc_hd__decap_3 PHY_724 ();
 sky130_fd_sc_hd__decap_3 PHY_725 ();
 sky130_fd_sc_hd__decap_3 PHY_726 ();
 sky130_fd_sc_hd__decap_3 PHY_727 ();
 sky130_fd_sc_hd__decap_3 PHY_728 ();
 sky130_fd_sc_hd__decap_3 PHY_729 ();
 sky130_fd_sc_hd__decap_3 PHY_730 ();
 sky130_fd_sc_hd__decap_3 PHY_731 ();
 sky130_fd_sc_hd__decap_3 PHY_732 ();
 sky130_fd_sc_hd__decap_3 PHY_733 ();
 sky130_fd_sc_hd__decap_3 PHY_734 ();
 sky130_fd_sc_hd__decap_3 PHY_735 ();
 sky130_fd_sc_hd__decap_3 PHY_736 ();
 sky130_fd_sc_hd__decap_3 PHY_737 ();
 sky130_fd_sc_hd__decap_3 PHY_738 ();
 sky130_fd_sc_hd__decap_3 PHY_739 ();
 sky130_fd_sc_hd__decap_3 PHY_740 ();
 sky130_fd_sc_hd__decap_3 PHY_741 ();
 sky130_fd_sc_hd__decap_3 PHY_742 ();
 sky130_fd_sc_hd__decap_3 PHY_743 ();
 sky130_fd_sc_hd__decap_3 PHY_744 ();
 sky130_fd_sc_hd__decap_3 PHY_745 ();
 sky130_fd_sc_hd__decap_3 PHY_746 ();
 sky130_fd_sc_hd__decap_3 PHY_747 ();
 sky130_fd_sc_hd__decap_3 PHY_748 ();
 sky130_fd_sc_hd__decap_3 PHY_749 ();
 sky130_fd_sc_hd__decap_3 PHY_750 ();
 sky130_fd_sc_hd__decap_3 PHY_751 ();
 sky130_fd_sc_hd__decap_3 PHY_752 ();
 sky130_fd_sc_hd__decap_3 PHY_753 ();
 sky130_fd_sc_hd__decap_3 PHY_754 ();
 sky130_fd_sc_hd__decap_3 PHY_755 ();
 sky130_fd_sc_hd__decap_3 PHY_756 ();
 sky130_fd_sc_hd__decap_3 PHY_757 ();
 sky130_fd_sc_hd__decap_3 PHY_758 ();
 sky130_fd_sc_hd__decap_3 PHY_759 ();
 sky130_fd_sc_hd__decap_3 PHY_760 ();
 sky130_fd_sc_hd__decap_3 PHY_761 ();
 sky130_fd_sc_hd__decap_3 PHY_762 ();
 sky130_fd_sc_hd__decap_3 PHY_763 ();
 sky130_fd_sc_hd__decap_3 PHY_764 ();
 sky130_fd_sc_hd__decap_3 PHY_765 ();
 sky130_fd_sc_hd__decap_3 PHY_766 ();
 sky130_fd_sc_hd__decap_3 PHY_767 ();
 sky130_fd_sc_hd__decap_3 PHY_768 ();
 sky130_fd_sc_hd__decap_3 PHY_769 ();
 sky130_fd_sc_hd__decap_3 PHY_770 ();
 sky130_fd_sc_hd__decap_3 PHY_771 ();
 sky130_fd_sc_hd__decap_3 PHY_772 ();
 sky130_fd_sc_hd__decap_3 PHY_773 ();
 sky130_fd_sc_hd__decap_3 PHY_774 ();
 sky130_fd_sc_hd__decap_3 PHY_775 ();
 sky130_fd_sc_hd__decap_3 PHY_776 ();
 sky130_fd_sc_hd__decap_3 PHY_777 ();
 sky130_fd_sc_hd__decap_3 PHY_778 ();
 sky130_fd_sc_hd__decap_3 PHY_779 ();
 sky130_fd_sc_hd__decap_3 PHY_780 ();
 sky130_fd_sc_hd__decap_3 PHY_781 ();
 sky130_fd_sc_hd__decap_3 PHY_782 ();
 sky130_fd_sc_hd__decap_3 PHY_783 ();
 sky130_fd_sc_hd__decap_3 PHY_784 ();
 sky130_fd_sc_hd__decap_3 PHY_785 ();
 sky130_fd_sc_hd__decap_3 PHY_786 ();
 sky130_fd_sc_hd__decap_3 PHY_787 ();
 sky130_fd_sc_hd__decap_3 PHY_788 ();
 sky130_fd_sc_hd__decap_3 PHY_789 ();
 sky130_fd_sc_hd__decap_3 PHY_790 ();
 sky130_fd_sc_hd__decap_3 PHY_791 ();
 sky130_fd_sc_hd__decap_3 PHY_792 ();
 sky130_fd_sc_hd__decap_3 PHY_793 ();
 sky130_fd_sc_hd__decap_3 PHY_794 ();
 sky130_fd_sc_hd__decap_3 PHY_795 ();
 sky130_fd_sc_hd__decap_3 PHY_796 ();
 sky130_fd_sc_hd__decap_3 PHY_797 ();
 sky130_fd_sc_hd__decap_3 PHY_798 ();
 sky130_fd_sc_hd__decap_3 PHY_799 ();
 sky130_fd_sc_hd__decap_3 PHY_800 ();
 sky130_fd_sc_hd__decap_3 PHY_801 ();
 sky130_fd_sc_hd__decap_3 PHY_802 ();
 sky130_fd_sc_hd__decap_3 PHY_803 ();
 sky130_fd_sc_hd__decap_3 PHY_804 ();
 sky130_fd_sc_hd__decap_3 PHY_805 ();
 sky130_fd_sc_hd__decap_3 PHY_806 ();
 sky130_fd_sc_hd__decap_3 PHY_807 ();
 sky130_fd_sc_hd__decap_3 PHY_808 ();
 sky130_fd_sc_hd__decap_3 PHY_809 ();
 sky130_fd_sc_hd__decap_3 PHY_810 ();
 sky130_fd_sc_hd__decap_3 PHY_811 ();
 sky130_fd_sc_hd__decap_3 PHY_812 ();
 sky130_fd_sc_hd__decap_3 PHY_813 ();
 sky130_fd_sc_hd__decap_3 PHY_814 ();
 sky130_fd_sc_hd__decap_3 PHY_815 ();
 sky130_fd_sc_hd__decap_3 PHY_816 ();
 sky130_fd_sc_hd__decap_3 PHY_817 ();
 sky130_fd_sc_hd__decap_3 PHY_818 ();
 sky130_fd_sc_hd__decap_3 PHY_819 ();
 sky130_fd_sc_hd__decap_3 PHY_820 ();
 sky130_fd_sc_hd__decap_3 PHY_821 ();
 sky130_fd_sc_hd__decap_3 PHY_822 ();
 sky130_fd_sc_hd__decap_3 PHY_823 ();
 sky130_fd_sc_hd__decap_3 PHY_824 ();
 sky130_fd_sc_hd__decap_3 PHY_825 ();
 sky130_fd_sc_hd__decap_3 PHY_826 ();
 sky130_fd_sc_hd__decap_3 PHY_827 ();
 sky130_fd_sc_hd__decap_3 PHY_828 ();
 sky130_fd_sc_hd__decap_3 PHY_829 ();
 sky130_fd_sc_hd__decap_3 PHY_830 ();
 sky130_fd_sc_hd__decap_3 PHY_831 ();
 sky130_fd_sc_hd__decap_3 PHY_832 ();
 sky130_fd_sc_hd__decap_3 PHY_833 ();
 sky130_fd_sc_hd__decap_3 PHY_834 ();
 sky130_fd_sc_hd__decap_3 PHY_835 ();
 sky130_fd_sc_hd__decap_3 PHY_836 ();
 sky130_fd_sc_hd__decap_3 PHY_837 ();
 sky130_fd_sc_hd__decap_3 PHY_838 ();
 sky130_fd_sc_hd__decap_3 PHY_839 ();
 sky130_fd_sc_hd__decap_3 PHY_840 ();
 sky130_fd_sc_hd__decap_3 PHY_841 ();
 sky130_fd_sc_hd__decap_3 PHY_842 ();
 sky130_fd_sc_hd__decap_3 PHY_843 ();
 sky130_fd_sc_hd__decap_3 PHY_844 ();
 sky130_fd_sc_hd__decap_3 PHY_845 ();
 sky130_fd_sc_hd__decap_3 PHY_846 ();
 sky130_fd_sc_hd__decap_3 PHY_847 ();
 sky130_fd_sc_hd__decap_3 PHY_848 ();
 sky130_fd_sc_hd__decap_3 PHY_849 ();
 sky130_fd_sc_hd__decap_3 PHY_850 ();
 sky130_fd_sc_hd__decap_3 PHY_851 ();
 sky130_fd_sc_hd__decap_3 PHY_852 ();
 sky130_fd_sc_hd__decap_3 PHY_853 ();
 sky130_fd_sc_hd__decap_3 PHY_854 ();
 sky130_fd_sc_hd__decap_3 PHY_855 ();
 sky130_fd_sc_hd__decap_3 PHY_856 ();
 sky130_fd_sc_hd__decap_3 PHY_857 ();
 sky130_fd_sc_hd__decap_3 PHY_858 ();
 sky130_fd_sc_hd__decap_3 PHY_859 ();
 sky130_fd_sc_hd__decap_3 PHY_860 ();
 sky130_fd_sc_hd__decap_3 PHY_861 ();
 sky130_fd_sc_hd__decap_3 PHY_862 ();
 sky130_fd_sc_hd__decap_3 PHY_863 ();
 sky130_fd_sc_hd__decap_3 PHY_864 ();
 sky130_fd_sc_hd__decap_3 PHY_865 ();
 sky130_fd_sc_hd__decap_3 PHY_866 ();
 sky130_fd_sc_hd__decap_3 PHY_867 ();
 sky130_fd_sc_hd__decap_3 PHY_868 ();
 sky130_fd_sc_hd__decap_3 PHY_869 ();
 sky130_fd_sc_hd__decap_3 PHY_870 ();
 sky130_fd_sc_hd__decap_3 PHY_871 ();
 sky130_fd_sc_hd__decap_3 PHY_872 ();
 sky130_fd_sc_hd__decap_3 PHY_873 ();
 sky130_fd_sc_hd__decap_3 PHY_874 ();
 sky130_fd_sc_hd__decap_3 PHY_875 ();
 sky130_fd_sc_hd__decap_3 PHY_876 ();
 sky130_fd_sc_hd__decap_3 PHY_877 ();
 sky130_fd_sc_hd__decap_3 PHY_878 ();
 sky130_fd_sc_hd__decap_3 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21432 ();
 sky130_fd_sc_hd__buf_12 input1 (.A(addr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_16 input2 (.A(addr[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_8 input3 (.A(data[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_16 input4 (.A(data[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(data[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(data[3]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(enb),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_16 input8 (.A(wr),
    .X(net8));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(r_data[0]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(r_data[1]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(r_data[2]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(r_data[3]));
 sky130_fd_sc_hd__conb_1 dff_ram_13 (.LO(net13));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_018_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_030_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\mem[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\mem[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\mem[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\mem[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net4));
 assign r_data[10] = net19;
 assign r_data[11] = net20;
 assign r_data[12] = net21;
 assign r_data[13] = net22;
 assign r_data[14] = net23;
 assign r_data[15] = net24;
 assign r_data[16] = net25;
 assign r_data[17] = net26;
 assign r_data[18] = net27;
 assign r_data[19] = net28;
 assign r_data[20] = net29;
 assign r_data[21] = net30;
 assign r_data[22] = net31;
 assign r_data[23] = net32;
 assign r_data[24] = net33;
 assign r_data[25] = net34;
 assign r_data[26] = net35;
 assign r_data[27] = net36;
 assign r_data[28] = net37;
 assign r_data[29] = net38;
 assign r_data[30] = net39;
 assign r_data[31] = net40;
 assign r_data[32] = net41;
 assign r_data[33] = net42;
 assign r_data[34] = net43;
 assign r_data[35] = net44;
 assign r_data[36] = net45;
 assign r_data[37] = net46;
 assign r_data[38] = net47;
 assign r_data[39] = net48;
 assign r_data[40] = net49;
 assign r_data[41] = net50;
 assign r_data[42] = net51;
 assign r_data[43] = net52;
 assign r_data[44] = net53;
 assign r_data[45] = net54;
 assign r_data[46] = net55;
 assign r_data[47] = net56;
 assign r_data[48] = net57;
 assign r_data[49] = net58;
 assign r_data[4] = net13;
 assign r_data[50] = net59;
 assign r_data[51] = net60;
 assign r_data[52] = net61;
 assign r_data[53] = net62;
 assign r_data[54] = net63;
 assign r_data[55] = net64;
 assign r_data[56] = net65;
 assign r_data[57] = net66;
 assign r_data[58] = net67;
 assign r_data[59] = net68;
 assign r_data[5] = net14;
 assign r_data[60] = net69;
 assign r_data[61] = net70;
 assign r_data[62] = net71;
 assign r_data[63] = net72;
 assign r_data[64] = net73;
 assign r_data[65] = net74;
 assign r_data[66] = net75;
 assign r_data[67] = net76;
 assign r_data[68] = net77;
 assign r_data[69] = net78;
 assign r_data[6] = net15;
 assign r_data[70] = net79;
 assign r_data[71] = net80;
 assign r_data[7] = net16;
 assign r_data[8] = net17;
 assign r_data[9] = net18;
endmodule
